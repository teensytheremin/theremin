* ADG752 SPICE Macro-model
* Generic Desc: CMOS, Low Voltage SPDT Switch
* Developed by: MPorley / ADGT
* Revision History: 1.0 (1/2018)
* Copyright 2018 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance of the terms and provisions in the License Statement.
*
* Begin Notes:
* The model will work on Vdd/Vss from 2.7V to 5.5V single supply.
* The model provides parametric specifications at +5V only and is not variable with Vdd. Please see datasheet page 3.
*
* Not Modeled:
*
* Parameters modeled include:
*	On Resistance
*	Ton and Toff
*	Break-Before-Make
*	Off Isolation
*	Crosstalk
*	Supply Currents: Iss/Idd
*	Bandwidth
*	Charge Injection
* Connections
*      1  = D1
*      2  = S1
*      3  = GND
*      4  = VDD
*      5  = NC
*      6  = IN1
*      8  = S2
*
.SUBCKT ADG752 5 8 3 6 5 2 4 1

.MODEL VON VSWITCH(Von=5 Voff=0.8 Ron=0.001 Roff=1000000000)
.MODEL VEN VSWITCH(Von=5 Voff=0.8 Ron=6000 Roff=7500)
.MODEL VNE VSWITCH(Von=5 Voff=0.8 Ron=16000 Roff=300)
.MODEL VRESET VSWITCH(Von=5 Voff=0.8 Ron=2700000 Roff=1000)
.MODEL DCLAMP D(IS=1E-15 IBV=1E-13)


* CROSSTALK
C12X 2 8 0.3E-012

* IDD/ISS
I1 4 3 0.001E-006

* Configuration: SPST 2:2


** SWITCH 1 **
*
* ESD PROTECTION DIODES
D11 3 1 DCLAMP
D12 1 4 DCLAMP
D13 3 2 DCLAMP
D14 2 4 DCLAMP
*
* OFF ISOLATION
C11 2 1 0.3E-012
*
* CHARGE INJECTION
C12 1 140 0.01E-012
C13 2 140 0.01E-012
*
* CD/CS OFF AND BANDWIDTH
C14 2 3 10E-012
C15 1 3 10e-012
*
* ON RESISTANCE
Ech155 1555 3 VALUE = { IF ((ABS(V(2)))>(ABS(V(184))),V(2),V(1)) }
R155 1555 3 1G
R11 137 1 0.001
S111 136 141 1141 3 VON
Ech111 1141 3 VALUE = { IF (V(1555)<1.3,5,0) }
Ech11 141 3 VALUE = { IF (V(1555)<1.3,0.294117647058824*(V(1555)-1.3)+10,0) }
S112 136 146 1146 3 VON
Ech112 1146 3 VALUE = { IF ((V(1555)>=1.3) & (V(1555)<=4),5,0) }
Ech12 146 3 VALUE = { IF ((V(1555)>=1.3) & (V(1555)<=4),((10-7)/((1.3-2.41837661840736)*(1.3-2.41837661840736)))*(V(1555)-2.41837661840736)*(V(1555)-2.41837661840736) + 7,0) }
S113 136 144 1144 3 VON
Ech113 1144 3 VALUE = { IF (V(1555)>4,5,0) }
Ech13 144 3 VALUE = { IF (V(1555)>4,-2*(V(1555)-4)+13,0) }
RIN1	136 3	1G
EOUT1 137 181	POLY(2) (136,3) (180,3) 0 0 0 0 0.999/1000
FCOPY1	3 180 VSENSE1 1
RSENSOR1 180 3	1K
VSENSE1 181 184	0
*
* TON/ TOFF/ BBM
S11 182 184 140 3 VON
S12 143 138 143 3 VEN
Ech14 143 3 VALUE = { IF(V(6)>=2.0, 5 , 0.8 ) }
eV1 140 3 138 3 1
C16 138 3 1e-012
*
* VOLTAGE SUPPLY REQUIREMENT
S13 2 182 185 3 VON
S15 139 185 139 3 VON
Ech16 139 3 VALUE = { IF((V(3)>=-0.5 & (V(4)<=5.5 & V(4)>=2.7)), 5 , 0.01 ) }


** SWITCH 2 **
*
* ESD PROTECTION DIODES
D21 3 9 DCLAMP
D22 9 4 DCLAMP
D23 3 8 DCLAMP
D24 8 4 DCLAMP
*
* OFF ISOLATION
C21 8 1 0.3E-012
*
* CHARGE INJECTION
C23 8 240 0.01E-012
*
* CD/CS OFF AND BANDWIDTH
C24 8 3 10E-012
*
* ON RESISTANCE
Ech255 2555 3 VALUE = { IF ((ABS(V(8)))>(ABS(V(284))),V(8),V(9)) }
R255 2555 3 1G
R21 237 1 0.001
S221 236 241 2241 3 VON
Ech221 2241 3 VALUE = { IF (V(2555)<1.3,5,0) }
Ech21 241 3 VALUE = { IF (V(2555)<1.3,0.294117647058824*(V(2555)-1.3)+10,0) }
S222 236 246 2246 3 VON
Ech222 2246 3 VALUE = { IF ((V(2555)>=1.3) & (V(2555)<=4),5,0) }
Ech22 246 3 VALUE = { IF ((V(2555)>=1.3) & (V(2555)<=4),((10-7)/((1.3-2.41837661840736)*(1.3-2.41837661840736)))*(V(2555)-2.41837661840736)*(V(2555)-2.41837661840736) + 7,0) }
S223 236 244 2244 3 VON
Ech223 2244 3 VALUE = { IF (V(2555)>4,5,0) }
Ech23 244 3 VALUE = { IF (V(2555)>4,-2*(V(2555)-4)+13,0) }
RIN2	236 3	1G
EOUT2 237 281	POLY(2) (236,3) (280,3) 0 0 0 0 0.999/1000
FCOPY2	3 280 VSENSE2 1
RSENSOR2 280 3	1K
VSENSE2 281 284	0
*
* TON/ TOFF/ BBM
S21 282 284 240 3 VON
S22 243 238 243 3 VNE
Ech24 243 3 VALUE = { IF(V(6)<2.0, 5 , 0.8 ) }
eV2 240 3 238 3 1
C26 238 3 1e-012
*
* VOLTAGE SUPPLY REQUIREMENT
S23 8 282 285 3 VON
S25 239 285 239 3 VON
Ech26 239 3 VALUE = { IF((V(3)>=-0.5 & (V(4)<=5.5 & V(4)>=2.7)), 5 , 0.01 ) }

.ENDS ADG752
